10 20 4
F 2 1 6
W 2 2 9
H 0 0 5 0
* 4 4 0
X 4 5 10
* 4 3 0
* 5 4 0
